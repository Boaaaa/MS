package CONSTANTS is
   	constant M_const   : integer := 4;	
	constant N_const   : integer := 4;	
	constant F_const   : integer := 4;
	constant word_size : integer := 4;
end CONSTANTS;
