package CONSTANTS is

   constant N_BIT   : integer := 4;	
   	
end CONSTANTS;
