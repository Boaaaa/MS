package CONSTANTS is

   constant N_BIT   : integer := 4;	
   constant N_Block   : integer := 8;	
   	
end CONSTANTS;
