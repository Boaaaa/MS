package CONSTANTS is

   constant ALL_BITS   : integer := 32;	
  
   constant N_subdiv  : integer := 4;	
   	
end CONSTANTS;
