package CONSTANTS is

    constant A_BIT   : integer := 16;	
    constant B_BIT   : integer := 8;
    --constant F_BIT   : integer := B_BIT + A_BIT; --final bit

 end CONSTANTS;
 